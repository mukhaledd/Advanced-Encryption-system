library verilog;
use verilog.vl_types.all;
entity mixColumns_tb is
end mixColumns_tb;
