library verilog;
use verilog.vl_types.all;
entity KeyExpansion_tb is
end KeyExpansion_tb;
