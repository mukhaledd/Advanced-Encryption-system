library verilog;
use verilog.vl_types.all;
entity AES_Encrypt_t is
end AES_Encrypt_t;
