
module S_Box(
input [7:0] State,
output reg[7:0] SubState
);

always@(State)
 case (State)
      	   8'h00: SubState=8'h63;
	   8'h01: SubState=8'h7c;
	   8'h02: SubState=8'h77;
	   8'h03: SubState=8'h7b;
	   8'h04: SubState=8'hf2;
	   8'h05: SubState=8'h6b;
	   8'h06: SubState=8'h6f;
	   8'h07: SubState=8'hc5;
	   8'h08: SubState=8'h30;
	   8'h09: SubState=8'h01;
	   8'h0a: SubState=8'h67;
	   8'h0b: SubState=8'h2b;
	   8'h0c: SubState=8'hfe;
	   8'h0d: SubState=8'hd7;
	   8'h0e: SubState=8'hab;
	   8'h0f: SubState=8'h76;
	   8'h10: SubState=8'hca;
	   8'h11: SubState=8'h82;
	   8'h12: SubState=8'hc9;
	   8'h13: SubState=8'h7d;
	   8'h14: SubState=8'hfa;
	   8'h15: SubState=8'h59;
	   8'h16: SubState=8'h47;
	   8'h17: SubState=8'hf0;
	   8'h18: SubState=8'had;
	   8'h19: SubState=8'hd4;
	   8'h1a: SubState=8'ha2;
	   8'h1b: SubState=8'haf;
	   8'h1c: SubState=8'h9c;
	   8'h1d: SubState=8'ha4;
	   8'h1e: SubState=8'h72;
	   8'h1f: SubState=8'hc0;
	   8'h20: SubState=8'hb7;
	   8'h21: SubState=8'hfd;
	   8'h22: SubState=8'h93;
	   8'h23: SubState=8'h26;
	   8'h24: SubState=8'h36;
	   8'h25: SubState=8'h3f;
	   8'h26: SubState=8'hf7;
	   8'h27: SubState=8'hcc;
	   8'h28: SubState=8'h34;
	   8'h29: SubState=8'ha5;
	   8'h2a: SubState=8'he5;
	   8'h2b: SubState=8'hf1;
	   8'h2c: SubState=8'h71;
	   8'h2d: SubState=8'hd8;
	   8'h2e: SubState=8'h31;
	   8'h2f: SubState=8'h15;
	   8'h30: SubState=8'h04;
	   8'h31: SubState=8'hc7;
	   8'h32: SubState=8'h23;
	   8'h33: SubState=8'hc3;
	   8'h34: SubState=8'h18;
	   8'h35: SubState=8'h96;
	   8'h36: SubState=8'h05;
	   8'h37: SubState=8'h9a;
	   8'h38: SubState=8'h07;
	   8'h39: SubState=8'h12;
	   8'h3a: SubState=8'h80;
	   8'h3b: SubState=8'he2;
	   8'h3c: SubState=8'heb;
	   8'h3d: SubState=8'h27;
	   8'h3e: SubState=8'hb2;
	   8'h3f: SubState=8'h75;
	   8'h40: SubState=8'h09;
	   8'h41: SubState=8'h83;
	   8'h42: SubState=8'h2c;
	   8'h43: SubState=8'h1a;
	   8'h44: SubState=8'h1b;
	   8'h45: SubState=8'h6e;
	   8'h46: SubState=8'h5a;
	   8'h47: SubState=8'ha0;
	   8'h48: SubState=8'h52;
	   8'h49: SubState=8'h3b;
	   8'h4a: SubState=8'hd6;
	   8'h4b: SubState=8'hb3;
	   8'h4c: SubState=8'h29;
	   8'h4d: SubState=8'he3;
	   8'h4e: SubState=8'h2f;
	   8'h4f: SubState=8'h84;
	   8'h50: SubState=8'h53;
	   8'h51: SubState=8'hd1;
	   8'h52: SubState=8'h00;
	   8'h53: SubState=8'hed;
	   8'h54: SubState=8'h20;
	   8'h55: SubState=8'hfc;
	   8'h56: SubState=8'hb1;
	   8'h57: SubState=8'h5b;
	   8'h58: SubState=8'h6a;
	   8'h59: SubState=8'hcb;
	   8'h5a: SubState=8'hbe;
	   8'h5b: SubState=8'h39;
	   8'h5c: SubState=8'h4a;
	   8'h5d: SubState=8'h4c;
	   8'h5e: SubState=8'h58;
	   8'h5f: SubState=8'hcf;
	   8'h60: SubState=8'hd0;
	   8'h61: SubState=8'hef;
	   8'h62: SubState=8'haa;
	   8'h63: SubState=8'hfb;
	   8'h64: SubState=8'h43;
	   8'h65: SubState=8'h4d;
	   8'h66: SubState=8'h33;
	   8'h67: SubState=8'h85;
	   8'h68: SubState=8'h45;
	   8'h69: SubState=8'hf9;
	   8'h6a: SubState=8'h02;
	   8'h6b: SubState=8'h7f;
	   8'h6c: SubState=8'h50;
	   8'h6d: SubState=8'h3c;
	   8'h6e: SubState=8'h9f;
	   8'h6f: SubState=8'ha8;
	   8'h70: SubState=8'h51;
	   8'h71: SubState=8'ha3;
	   8'h72: SubState=8'h40;
	   8'h73: SubState=8'h8f;
	   8'h74: SubState=8'h92;
	   8'h75: SubState=8'h9d;
	   8'h76: SubState=8'h38;
	   8'h77: SubState=8'hf5;
	   8'h78: SubState=8'hbc;
	   8'h79: SubState=8'hb6;
	   8'h7a: SubState=8'hda;
	   8'h7b: SubState=8'h21;
	   8'h7c: SubState=8'h10;
	   8'h7d: SubState=8'hff;
	   8'h7e: SubState=8'hf3;
	   8'h7f: SubState=8'hd2;
	   8'h80: SubState=8'hcd;
	   8'h81: SubState=8'h0c;
	   8'h82: SubState=8'h13;
	   8'h83: SubState=8'hec;
	   8'h84: SubState=8'h5f;
	   8'h85: SubState=8'h97;
	   8'h86: SubState=8'h44;
	   8'h87: SubState=8'h17;
	   8'h88: SubState=8'hc4;
	   8'h89: SubState=8'ha7;
	   8'h8a: SubState=8'h7e;
	   8'h8b: SubState=8'h3d;
	   8'h8c: SubState=8'h64;
	   8'h8d: SubState=8'h5d;
	   8'h8e: SubState=8'h19;
	   8'h8f: SubState=8'h73;
	   8'h90: SubState=8'h60;
	   8'h91: SubState=8'h81;
	   8'h92: SubState=8'h4f;
	   8'h93: SubState=8'hdc;
	   8'h94: SubState=8'h22;
	   8'h95: SubState=8'h2a;
	   8'h96: SubState=8'h90;
	   8'h97: SubState=8'h88;
	   8'h98: SubState=8'h46;
	   8'h99: SubState=8'hee;
	   8'h9a: SubState=8'hb8;
	   8'h9b: SubState=8'h14;
	   8'h9c: SubState=8'hde;
	   8'h9d: SubState=8'h5e;
	   8'h9e: SubState=8'h0b;
	   8'h9f: SubState=8'hdb;
	   8'ha0: SubState=8'he0;
	   8'ha1: SubState=8'h32;
	   8'ha2: SubState=8'h3a;
	   8'ha3: SubState=8'h0a;
	   8'ha4: SubState=8'h49;
	   8'ha5: SubState=8'h06;
	   8'ha6: SubState=8'h24;
	   8'ha7: SubState=8'h5c;
	   8'ha8: SubState=8'hc2;
	   8'ha9: SubState=8'hd3;
	   8'haa: SubState=8'hac;
	   8'hab: SubState=8'h62;
	   8'hac: SubState=8'h91;
	   8'had: SubState=8'h95;
	   8'hae: SubState=8'he4;
	   8'haf: SubState=8'h79;
	   8'hb0: SubState=8'he7;
	   8'hb1: SubState=8'hc8;
	   8'hb2: SubState=8'h37;
	   8'hb3: SubState=8'h6d;
	   8'hb4: SubState=8'h8d;
	   8'hb5: SubState=8'hd5;
	   8'hb6: SubState=8'h4e;
	   8'hb7: SubState=8'ha9;
	   8'hb8: SubState=8'h6c;
	   8'hb9: SubState=8'h56;
	   8'hba: SubState=8'hf4;
	   8'hbb: SubState=8'hea;
	   8'hbc: SubState=8'h65;
	   8'hbd: SubState=8'h7a;
	   8'hbe: SubState=8'hae;
	   8'hbf: SubState=8'h08;
	   8'hc0: SubState=8'hba;
	   8'hc1: SubState=8'h78;
	   8'hc2: SubState=8'h25;
	   8'hc3: SubState=8'h2e;
	   8'hc4: SubState=8'h1c;
	   8'hc5: SubState=8'ha6;
	   8'hc6: SubState=8'hb4;
	   8'hc7: SubState=8'hc6;
	   8'hc8: SubState=8'he8;
	   8'hc9: SubState=8'hdd;
	   8'hca: SubState=8'h74;
	   8'hcb: SubState=8'h1f;
	   8'hcc: SubState=8'h4b;
	   8'hcd: SubState=8'hbd;
	   8'hce: SubState=8'h8b;
	   8'hcf: SubState=8'h8a;
	   8'hd0: SubState=8'h70;
	   8'hd1: SubState=8'h3e;
	   8'hd2: SubState=8'hb5;
	   8'hd3: SubState=8'h66;
	   8'hd4: SubState=8'h48;
	   8'hd5: SubState=8'h03;
	   8'hd6: SubState=8'hf6;
	   8'hd7: SubState=8'h0e;
	   8'hd8: SubState=8'h61;
	   8'hd9: SubState=8'h35;
	   8'hda: SubState=8'h57;
	   8'hdb: SubState=8'hb9;
	   8'hdc: SubState=8'h86;
	   8'hdd: SubState=8'hc1;
	   8'hde: SubState=8'h1d;
	   8'hdf: SubState=8'h9e;
	   8'he0: SubState=8'he1;
	   8'he1: SubState=8'hf8;
	   8'he2: SubState=8'h98;
	   8'he3: SubState=8'h11;
	   8'he4: SubState=8'h69;
	   8'he5: SubState=8'hd9;
	   8'he6: SubState=8'h8e;
	   8'he7: SubState=8'h94;
	   8'he8: SubState=8'h9b;
	   8'he9: SubState=8'h1e;
	   8'hea: SubState=8'h87;
	   8'heb: SubState=8'he9;
	   8'hec: SubState=8'hce;
	   8'hed: SubState=8'h55;
	   8'hee: SubState=8'h28;
	   8'hef: SubState=8'hdf;
	   8'hf0: SubState=8'h8c;
	   8'hf1: SubState=8'ha1;
	   8'hf2: SubState=8'h89;
	   8'hf3: SubState=8'h0d;
	   8'hf4: SubState=8'hbf;
	   8'hf5: SubState=8'he6;
	   8'hf6: SubState=8'h42;
	   8'hf7: SubState=8'h68;
	   8'hf8: SubState=8'h41;
	   8'hf9: SubState=8'h99;
	   8'hfa: SubState=8'h2d;
	   8'hfb: SubState=8'h0f;
	   8'hfc: SubState=8'hb0;
	   8'hfd: SubState=8'h54;
	   8'hfe: SubState=8'hbb;
	   8'hff: SubState=8'h16;
	endcase

endmodule