library verilog;
use verilog.vl_types.all;
entity Add_Round_Key_tb is
end Add_Round_Key_tb;
