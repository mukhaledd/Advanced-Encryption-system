library verilog;
use verilog.vl_types.all;
entity AES_Encryption_tb is
end AES_Encryption_tb;
