library verilog;
use verilog.vl_types.all;
entity ShiftRows_tb is
end ShiftRows_tb;
