library verilog;
use verilog.vl_types.all;
entity Sub_Bytes_tb is
end Sub_Bytes_tb;
